`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:35:03 04/10/2017 
// Design Name: 
// Module Name:    SSEGDriver 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SSEGDriver(input clk,
						input [7:0] digit1,
						input [7:0] digit2,
						input [7:0] digit3,
						input [7:0] digit4,
						output reg [3:0] SSEGD,
						output reg [7:0] SSEG);


endmodule
